module geometry
